module InputFeeder(

	output reg [6:0] out,
	input clk

	);
	
	integer address_pointer;
	
	reg [6:0] InputBuffer [0:5];
	
	initial begin
	
		address_pointer <= 0;
		
		out <= 7'b1111111;
		
		$readmemb("Fifo_Input.txt", InputBuffer);
		
	end
	
	always @(posedge clk) begin
	
		if (address_pointer < 6) begin
		
			out <= InputBuffer[address_pointer];
			
			address_pointer = address_pointer + 1;
			
		end else begin
		
			address_pointer = 0;
			
		end
		
	end
	
endmodule

//=======================================================
//  This code is generated by Terasic System Builder
//=======================================================

module Lab1_Part3(

	//////////// ADC //////////
	output		          		ADC_CONVST,
	output		          		ADC_DIN,
	input 		          		ADC_DOUT,
	output		          		ADC_SCLK,

	//////////// Audio //////////
	input 		          		AUD_ADCDAT,
	inout 		          		AUD_ADCLRCK,
	inout 		          		AUD_BCLK,
	output		          		AUD_DACDAT,
	inout 		          		AUD_DACLRCK,
	output		          		AUD_XCK,

	//////////// CLOCK //////////
	input 		          		CLOCK2_50,
	input 		          		CLOCK3_50,
	input 		          		CLOCK4_50,
	input 		          		CLOCK_50,

	//////////// SDRAM //////////
	output		    [12:0]		DRAM_ADDR,
	output		     [1:0]		DRAM_BA,
	output		          		DRAM_CAS_N,
	output		          		DRAM_CKE,
	output		          		DRAM_CLK,
	output		          		DRAM_CS_N,
	inout 		    [15:0]		DRAM_DQ,
	output		          		DRAM_LDQM,
	output		          		DRAM_RAS_N,
	output		          		DRAM_UDQM,
	output		          		DRAM_WE_N,

	//////////// I2C for Audio and Video-In //////////
	output		          		FPGA_I2C_SCLK,
	inout 		          		FPGA_I2C_SDAT,

	//////////// SEG7 //////////
	output		     [6:0]		HEX0,
	output		     [6:0]		HEX1,
	output		     [6:0]		HEX2,
	output		     [6:0]		HEX3,
	output		     [6:0]		HEX4,
	output		     [6:0]		HEX5,

	//////////// IR //////////
	input 		          		IRDA_RXD,
	output		          		IRDA_TXD,

	//////////// KEY //////////
	input 		     [3:0]		KEY,

	//////////// LED //////////
	output		     [9:0]		LEDR,

	//////////// PS2 //////////
	inout 		          		PS2_CLK,
	inout 		          		PS2_CLK2,
	inout 		          		PS2_DAT,
	inout 		          		PS2_DAT2,

	//////////// SW //////////
	input 		     [9:0]		SW,

	//////////// Video-In //////////
	input 		          		TD_CLK27,
	input 		     [7:0]		TD_DATA,
	input 		          		TD_HS,
	output		          		TD_RESET_N,
	input 		          		TD_VS,

	//////////// VGA //////////
	output		          		VGA_BLANK_N,
	output		     [7:0]		VGA_B,
	output		          		VGA_CLK,
	output		     [7:0]		VGA_G,
	output		          		VGA_HS,
	output		     [7:0]		VGA_R,
	output		          		VGA_SYNC_N,
	output		          		VGA_VS
);



//=======================================================
//  REG/WIRE declarations
//=======================================================

	reg [6:0] hex0_buffer, hex1_buffer, hex2_buffer, hex3_buffer, hex4_buffer, hex5_buffer;
	reg [9:0] sw_buffer;
	reg clk_slow, clk_fast;
	reg [24:0] counter, counter1;
	
	wire [6:0] out;
	wire current_clk;

//=======================================================
//  Structural coding
//=======================================================

/*

	To-do:
	
	1) One push button will reset the entire system.
	2) One push button will invert the patterns on both the LEDs and the 7-segment displays (on → off, off → on)
	3) One push button will speed up the horizontal scrolling movement displayed on the seven segment display. You choose how fast
	4) One push button will pause the horizontal scrolling movement displayed on the seven segment display. Pushing the pause again will continue the scrolling movement. 
		While in the pause state, other push buttons will have no effect on the seven segment display behavior. However, the user can still use the switches to change the red LED
		pattern at anytime.

*/

	//clk_slow divider-1Hz 

	always @(posedge CLOCK_50) begin

		if (counter == 24999999) begin
		
			counter <= 0;
			
			clk_slow <= ~clk_slow;
			
		end else begin
		
			counter <= counter + 1;
			
		end
		
	end

	//clk_fast divider-5Hz 

	always @(posedge CLOCK_50) begin

		if (counter1 == 9999999) begin
		
			counter1 <= 0;
			
			clk_fast <= ~clk_fast;
			
		end else begin
		
			counter1 <= counter1 + 1;
			
		end
		
	end
	
	InputFeeder u0 (.clk(current_clk), .out(out));
	
	assign current_clk = (KEY[1] == 0) ? clk_fast : clk_slow; //use KEY1 to choose between clock speeds, so we can speed up the display

	always @(posedge current_clk) begin
		
		if (KEY[3] == 0) begin //reset
		
			hex0_buffer <= 7'b1111111;
			hex1_buffer <= 7'b1111111;
			hex2_buffer <= 7'b1111111;
			hex3_buffer <= 7'b1111111;
			hex4_buffer <= 7'b1111111;
			hex5_buffer <= 7'b1111111;
		
		end
		
		else if (KEY[2] == 0) begin //invert switch and displays
		
			sw_buffer <= ~SW;
			
			hex5_buffer <= out;
			hex4_buffer <= hex5_buffer;
			hex3_buffer <= hex4_buffer;
			hex2_buffer <= hex3_buffer;
			hex1_buffer <= hex2_buffer;
			hex0_buffer <= hex1_buffer;
		
		end
		
		else if (KEY[0] == 0) begin //pause everything
		
			hex5_buffer <= hex5_buffer;
			hex4_buffer <= hex4_buffer;
			hex3_buffer <= hex3_buffer;
			hex2_buffer <= hex2_buffer;
			hex1_buffer <= hex1_buffer;
			hex0_buffer <= hex0_buffer;
			
			sw_buffer <= SW;
		
		end
			
		else begin
		
			//default case
			hex0_buffer <= out;
			hex1_buffer <= hex0_buffer;
			hex2_buffer <= hex1_buffer;
			hex3_buffer <= hex2_buffer;
			hex4_buffer <= hex3_buffer;
			hex5_buffer <= hex4_buffer;
			
			sw_buffer <= SW;
			
		end
		
	end
	
	assign HEX0 = hex0_buffer;
	assign HEX1 = hex1_buffer;
	assign HEX2 = hex2_buffer;
	assign HEX3 = hex3_buffer;
	assign HEX4 = hex4_buffer;
	assign HEX5 = hex5_buffer;
	
	assign LEDR = sw_buffer;

endmodule
