module InputFeeder(

	output reg [6:0] out,
	input clk
	
); 

	reg [6:0] inputBuffer [0:5]; //6 lines of 7 bits each
	
	integer address_pointer;
	
	initial begin 
		
		$readmemb("FIFO_Input.txt", inputBuffer);
		
		address_pointer = 0;
		
		out = 7'b1111111;
		
	end

	always @(posedge clk) begin	

		if (address_pointer < 6) begin
		
		out <= inputBuffer[address_pointer];
		
		address_pointer <= address_pointer + 1;
		
		end else begin
		
		address_pointer = 0;
		
		end
		
	end
	
endmodule

//=======================================================
//  This code is generated by Terasic System Builder
//=======================================================

module Lab1_Part2(

	//////////// ADC //////////
	output		          		ADC_CONVST,
	output		          		ADC_DIN,
	input 		          		ADC_Dout,
	output		          		ADC_SCLK,

	//////////// Audio //////////
	input 		          		AUD_ADCDAT,
	inout 		          		AUD_ADCLRCK,
	inout 		          		AUD_BCLK,
	output		          		AUD_DACDAT,
	inout 		          		AUD_DACLRCK,
	output		          		AUD_XCK,

	//////////// CLOCK //////////
	input 		          		CLOCK2_50,
	input 		          		CLOCK3_50,
	input 		          		CLOCK4_50,
	input 		          		CLOCK_50,

	//////////// SDRAM //////////
	output		    [12:0]		DRAM_ADDR,
	output		     [1:0]		DRAM_BA,
	output		          		DRAM_CAS_N,
	output		          		DRAM_CKE,
	output		          		DRAM_CLK,
	output		          		DRAM_CS_N,
	inout 		    [15:0]		DRAM_DQ,
	output		          		DRAM_LDQM,
	output		          		DRAM_RAS_N,
	output		          		DRAM_UDQM,
	output		          		DRAM_WE_N,

	//////////// I2C for Audio and Video-In //////////
	output		          		FPGA_I2C_SCLK,
	inout 		          		FPGA_I2C_SDAT,

	//////////// SEG7 //////////
	output		     [6:0]		HEX0,
	output		     [6:0]		HEX1,
	output		     [6:0]		HEX2,
	output		     [6:0]		HEX3,
	output		     [6:0]		HEX4,
	output		     [6:0]		HEX5,

	//////////// IR //////////
	input 		          		IRDA_RXD,
	output		          		IRDA_TXD,

	//////////// KEY //////////
	input 		     [3:0]		KEY,

	//////////// LED //////////
	output		     [9:0]		LEDR,

	//////////// PS2 //////////
	inout 		          		PS2_CLK,
	inout 		          		PS2_CLK2,
	inout 		          		PS2_DAT,
	inout 		          		PS2_DAT2,

	//////////// SW //////////
	input 		     [9:0]		SW,

	//////////// Video-In //////////
	input 		          		TD_CLK27,
	input 		     [7:0]		TD_DATA,
	input 		          		TD_HS,
	output		          		TD_RESET_N,
	input 		          		TD_VS,

	//////////// VGA //////////
	output		          		VGA_BLANK_N,
	output		     [7:0]		VGA_B,
	output		          		VGA_CLK,
	output		     [7:0]		VGA_G,
	output		          		VGA_HS,
	output		     [7:0]		VGA_R,
	output		          		VGA_SYNC_N,
	output		          		VGA_VS
);



//=======================================================
//  REG/WIRE declarations
//=======================================================

	reg [6:0] hex0_reg, hex1_reg, hex2_reg, hex3_reg, hex4_reg, hex5_reg;
	wire [6:0] out;
	reg [24:0] counter;
	reg slow_clk;

//=======================================================
//  Structural coding
//=======================================================
	
//  Clock divider for 1Hz

	always @(posedge CLOCK_50) begin
	
		if (counter == 24999999) begin
		
			counter <= 0;
			slow_clk <= ~slow_clk;
			
		end else begin
		
			counter <= counter + 1;
			
		end
		
	end
	
	InputFeeder u0(.out(out), .clk(slow_clk));
	
	always @(posedge slow_clk) begin
	
		hex5_reg <= hex4_reg;
		hex4_reg <= hex3_reg;
		hex3_reg <= hex2_reg;
		hex2_reg <= hex1_reg;
		hex1_reg <= hex0_reg;
		hex0_reg <= out;

end

		assign HEX0 = hex0_reg;
		assign HEX1 = hex1_reg;
		assign HEX2 = hex2_reg;
		assign HEX3 = hex3_reg;
		assign HEX4 = hex4_reg;
		assign HEX5 = hex5_reg;

endmodule
